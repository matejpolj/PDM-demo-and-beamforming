----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 26.07.2024 14:01:29
-- Design Name: 
-- Module Name: beam_gen - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package pkg is
    constant x_res : integer := 80;
    constant y_res : integer := 60;

    type delay_array    is array (natural range <>) of integer range 0 to 25;
    type delay_matrix   is array (natural range <>) of delay_array(0 to y_res-1);
    
    constant delay_matrix_1 : delay_matrix(0 to x_res-1) := ((25,24,24,24,24,23,23,23,23,22,22,22,22,22,22,21,21,21,21,21,21,21,21,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,21,21,21,21,21,21,21,22,22,22,22,22,22,23,23,23,23,24,24,24,24),
            (24,24,24,23,23,23,23,22,22,22,22,22,21,21,21,21,21,21,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,21,21,21,21,21,22,22,22,22,22,23,23,23,23,24,24),
            (24,23,23,23,23,22,22,22,22,21,21,21,21,21,21,20,20,20,20,20,20,20,20,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,20,20,20,20,20,20,20,20,21,21,21,21,21,21,22,22,22,22,23,23,23,23),
            (23,23,23,22,22,22,22,21,21,21,21,21,20,20,20,20,20,20,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,20,20,20,20,20,20,21,21,21,21,21,22,22,22,22,23,23),
            (23,22,22,22,22,21,21,21,21,20,20,20,20,20,20,19,19,19,19,19,19,19,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,19,19,19,19,19,19,19,20,20,20,20,20,20,21,21,21,21,22,22,22,22),
            (22,22,22,21,21,21,21,20,20,20,20,20,19,19,19,19,19,19,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,19,19,19,19,19,19,20,20,20,20,20,21,21,21,21,22,22),
            (22,22,21,21,21,20,20,20,20,20,19,19,19,19,19,18,18,18,18,18,18,18,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,18,18,18,18,18,18,18,19,19,19,19,19,20,20,20,20,20,21,21,21,22),
            (21,21,21,21,20,20,20,20,19,19,19,19,18,18,18,18,18,18,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,18,18,18,18,18,18,19,19,19,19,20,20,20,20,21,21,21),
            (21,21,20,20,20,20,19,19,19,19,18,18,18,18,18,17,17,17,17,17,17,17,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,17,17,17,17,17,17,18,18,18,18,18,19,19,19,19,20,20,20,20,21),
            (21,20,20,20,19,19,19,19,18,18,18,18,17,17,17,17,17,17,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,17,17,17,17,17,18,18,18,18,19,19,19,19,20,20,20),
            (20,20,19,19,19,19,18,18,18,18,17,17,17,17,17,16,16,16,16,16,16,16,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,17,17,17,17,17,18,18,18,18,19,19,19,19,20),
            (20,19,19,19,18,18,18,18,17,17,17,17,16,16,16,16,16,16,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,17,17,17,17,18,18,18,18,19,19,19),
            (19,19,19,18,18,18,17,17,17,17,16,16,16,16,16,15,15,15,15,15,15,15,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,16,16,16,16,16,17,17,17,17,18,18,18,19,19),
            (19,19,18,18,18,17,17,17,17,16,16,16,16,15,15,15,15,15,14,14,14,14,14,14,14,14,14,14,14,14,13,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,16,16,16,16,17,17,17,17,18,18,18,19),
            (18,18,18,17,17,17,17,16,16,16,16,15,15,15,15,14,14,14,14,14,14,14,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,15,15,15,15,16,16,16,16,17,17,17,17,18,18),
            (18,18,17,17,17,16,16,16,16,15,15,15,15,14,14,14,14,14,13,13,13,13,13,13,13,13,13,13,13,13,12,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,15,15,15,15,16,16,16,16,17,17,17,18),
            (18,17,17,17,16,16,16,15,15,15,15,14,14,14,14,14,13,13,13,13,13,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,14,14,14,14,14,15,15,15,15,16,16,16,17,17,17),
            (17,17,17,16,16,16,15,15,15,14,14,14,14,13,13,13,13,13,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,14,14,14,14,15,15,15,16,16,16,17,17),
            (17,17,16,16,16,15,15,15,14,14,14,14,13,13,13,13,12,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,13,13,13,13,14,14,14,14,15,15,15,16,16,16,17),
            (16,16,16,15,15,15,14,14,14,14,13,13,13,13,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,13,13,13,13,14,14,14,14,15,15,15,16,16),
            (16,16,15,15,15,14,14,14,13,13,13,13,12,12,12,12,12,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,12,12,12,12,12,13,13,13,13,14,14,14,15,15,15,16),
            (16,15,15,15,14,14,14,13,13,13,13,12,12,12,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,12,12,12,13,13,13,13,14,14,14,15,15,15),
            (15,15,15,14,14,14,13,13,13,12,12,12,12,11,11,11,11,10,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,11,11,11,11,12,12,12,12,13,13,13,14,14,14,15,15),
            (15,15,14,14,14,13,13,13,12,12,12,11,11,11,11,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,11,11,11,11,12,12,12,13,13,13,14,14,14,15),
            (15,14,14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,10,9,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,10,10,10,10,10,11,11,11,12,12,12,13,13,13,14,14,14),
            (14,14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,10,10,10,10,11,11,11,12,12,12,13,13,13,14,14),
            (14,14,13,13,13,12,12,11,11,11,11,10,10,10,9,9,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,9,9,9,9,9,10,10,10,11,11,11,11,12,12,13,13,13,14),
            (14,13,13,13,12,12,11,11,11,10,10,10,10,9,9,9,9,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,9,9,9,9,10,10,10,10,11,11,11,12,12,13,13,13),
            (13,13,13,12,12,11,11,11,10,10,10,9,9,9,9,8,8,8,8,7,7,7,7,7,7,7,7,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,8,8,8,8,9,9,9,9,10,10,10,11,11,11,12,12,13,13),
            (13,13,12,12,12,11,11,10,10,10,9,9,9,9,8,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,8,9,9,9,9,10,10,10,11,11,12,12,12,13),
            (13,12,12,12,11,11,10,10,10,9,9,9,8,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,12,12,12),
            (12,12,12,11,11,11,10,10,9,9,9,8,8,8,8,7,7,7,7,6,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,11,11,11,12,12),
            (12,12,11,11,11,10,10,9,9,9,8,8,8,7,7,7,7,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12),
            (12,12,11,11,10,10,10,9,9,8,8,8,7,7,7,7,6,6,6,6,5,5,5,5,5,5,5,4,4,4,4,4,4,4,5,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,10,10,10,11,11,12),
            (12,11,11,10,10,10,9,9,9,8,8,7,7,7,7,6,6,6,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,6,6,6,7,7,7,7,8,8,9,9,9,10,10,10,11,11),
            (11,11,11,10,10,9,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11),
            (11,11,10,10,10,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,4,4,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,10,11),
            (11,11,10,10,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,11),
            (11,10,10,10,9,9,8,8,7,7,7,6,6,6,5,5,5,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,10,10,10),
            (11,10,10,9,9,8,8,8,7,7,7,6,6,5,5,5,5,4,4,4,3,3,3,3,3,3,3,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,5,5,5,5,6,6,7,7,7,8,8,8,9,9,10,10),
            (10,10,10,9,9,8,8,7,7,7,6,6,6,5,5,5,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,10,10),
            (10,10,9,9,9,8,8,7,7,6,6,6,5,5,5,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,9,9,9,10),
            (10,10,9,9,8,8,8,7,7,6,6,6,5,5,4,4,4,4,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,4,4,4,4,5,5,6,6,6,7,7,8,8,8,9,9,10),
            (10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10),
            (10,9,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,9),
            (10,9,9,8,8,8,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,8,9,9),
            (10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (9,9,9,8,8,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,9,9),
            (9,9,9,8,8,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,9,9),
            (9,9,9,8,8,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,0,0,0,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,3,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,5,5,5,6,6,7,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9),
            (10,9,9,8,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,8,9,9),
            (10,10,9,9,8,8,7,7,6,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,9,9,10),
            (10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,2,2,1,1,1,1,1,2,2,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10),
            (10,10,9,9,8,8,8,7,7,6,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,8,9,9,10),
            (10,10,9,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,9,10),
            (11,10,10,9,9,8,8,8,7,7,6,6,6,5,5,5,4,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5,6,6,6,7,7,8,8,8,9,9,10,10),
            (11,10,10,9,9,9,8,8,7,7,7,6,6,6,5,5,5,4,4,4,4,3,3,3,3,3,3,3,3,3,2,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,9,10,10),
            (11,10,10,10,9,9,8,8,8,7,7,7,6,6,6,5,5,5,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,10),
            (11,11,10,10,9,9,9,8,8,7,7,7,6,6,6,6,5,5,5,4,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,6,6,6,6,7,7,7,8,8,9,9,9,10,10,11),
            (11,11,11,10,10,9,9,9,8,8,7,7,7,6,6,6,6,5,5,5,5,4,4,4,4,4,4,4,4,3,3,3,4,4,4,4,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,8,8,9,9,9,10,10,11,11),
            (12,11,11,10,10,10,9,9,8,8,8,7,7,7,6,6,6,6,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,8,8,8,9,9,10,10,10,11,11),
            (12,11,11,11,10,10,9,9,9,8,8,8,7,7,7,6,6,6,6,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,6,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11,11),
            (12,12,11,11,10,10,10,9,9,9,8,8,8,7,7,7,7,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,12),
            (12,12,12,11,11,10,10,10,9,9,9,8,8,8,7,7,7,7,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,12,12),
            (13,12,12,11,11,11,10,10,10,9,9,9,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,5,5,5,5,5,5,5,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12),
            (13,13,12,12,11,11,11,10,10,10,9,9,9,8,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13),
            (13,13,12,12,12,11,11,11,10,10,10,9,9,9,8,8,8,8,8,7,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,8,8,8,8,8,9,9,9,10,10,10,11,11,11,12,12,12,13),
            (14,13,13,12,12,12,11,11,11,10,10,10,9,9,9,9,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,9,9,9,9,10,10,10,11,11,11,12,12,12,13,13),
            (14,13,13,13,12,12,12,11,11,11,10,10,10,10,9,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,9,9,9,9,10,10,10,10,11,11,11,12,12,12,13,13,13),
            (14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,10,10,10,10,11,11,11,12,12,12,13,13,13,14),
            (15,14,14,13,13,13,12,12,12,11,11,11,11,10,10,10,10,9,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,10,10,10,10,11,11,11,11,12,12,12,13,13,13,14,14),
            (15,14,14,14,13,13,13,12,12,12,12,11,11,11,10,10,10,10,10,9,9,9,9,9,9,9,9,9,8,8,8,8,8,9,9,9,9,9,9,9,9,9,10,10,10,10,10,11,11,11,12,12,12,12,13,13,13,14,14,14));
    
    constant delay_matrix_2 : delay_matrix(0 to x_res-1) := ((17,16,16,16,16,16,15,15,15,15,15,15,15,15,15,15,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,17,17,17,17,18,18,18,18,19,19,19,20,20,20,21,21,21,22,22,22,23,23),
            (16,16,16,15,15,15,15,15,15,15,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,16,16,16,16,16,17,17,17,17,18,18,18,19,19,19,20,20,20,21,21,21,22,22,22,23),
            (16,15,15,15,15,15,14,14,14,14,14,14,14,14,14,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,16,16,16,16,17,17,17,18,18,18,19,19,19,19,20,20,21,21,21,22,22,22),
            (15,15,15,15,14,14,14,14,14,14,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,15,15,15,15,16,16,16,16,17,17,17,17,18,18,18,19,19,19,20,20,21,21,21,22,22),
            (15,14,14,14,14,14,14,13,13,13,13,13,13,13,13,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,14,14,14,14,14,15,15,15,15,16,16,16,16,17,17,17,18,18,18,19,19,19,20,20,21,21,21,22),
            (14,14,14,14,13,13,13,13,13,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,14,14,14,14,15,15,15,15,16,16,16,17,17,17,18,18,18,19,19,19,20,20,21,21,21),
            (14,14,13,13,13,13,13,12,12,12,12,12,12,12,12,12,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,13,13,13,13,13,14,14,14,14,15,15,15,16,16,16,17,17,17,18,18,18,19,19,19,20,20,21,21),
            (13,13,13,13,12,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,13,13,13,13,13,14,14,14,15,15,15,16,16,16,16,17,17,18,18,18,19,19,19,20,20,21),
            (13,13,12,12,12,12,12,11,11,11,11,11,11,11,11,11,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,12,12,12,12,12,13,13,13,13,14,14,14,14,15,15,15,16,16,16,17,17,18,18,18,19,19,20,20,20),
            (13,12,12,12,12,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,12,12,12,12,13,13,13,13,14,14,14,15,15,15,16,16,16,17,17,18,18,18,19,19,20,20),
            (12,12,12,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,9,9,9,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,12,12,12,12,13,13,13,14,14,14,15,15,15,16,16,16,17,17,18,18,18,19,19,20),
            (12,11,11,11,11,10,10,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,11,11,11,11,12,12,12,12,13,13,13,14,14,14,15,15,15,16,16,17,17,17,18,18,19,19,19),
            (11,11,11,11,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,11,11,11,11,12,12,12,13,13,13,14,14,14,15,15,15,16,16,17,17,17,18,18,19,19),
            (11,11,10,10,10,10,9,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,10,10,10,10,10,11,11,11,12,12,12,13,13,13,14,14,14,15,15,15,16,16,17,17,17,18,18,19),
            (10,10,10,10,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,10,10,10,10,11,11,11,12,12,12,13,13,13,14,14,14,15,15,16,16,16,17,17,18,18,18),
            (10,10,10,9,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,9,9,9,9,10,10,10,11,11,11,11,12,12,13,13,13,14,14,14,15,15,16,16,16,17,17,18,18),
            (10,9,9,9,9,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,9,9,9,10,10,10,10,11,11,11,12,12,13,13,13,14,14,14,15,15,16,16,17,17,17,18),
            (9,9,9,9,8,8,8,8,7,7,7,7,7,7,7,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,8,8,8,8,9,9,9,9,10,10,10,11,11,11,12,12,13,13,13,14,14,15,15,15,16,16,17,17,18),
            (9,9,8,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,8,8,8,9,9,9,9,10,10,10,11,11,12,12,12,13,13,13,14,14,15,15,16,16,17,17,17),
            (9,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,5,5,5,6,6,6,6,6,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,12,12,12,13,13,14,14,14,15,15,16,16,17,17),
            (8,8,8,7,7,7,7,6,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,13,14,14,15,15,16,16,16,17),
            (8,8,7,7,7,7,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,14,14,14,15,15,16,16,17),
            (8,7,7,7,6,6,6,6,5,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,10,10,10,11,11,12,12,12,13,13,14,14,15,15,16,16,16),
            (7,7,7,6,6,6,6,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,6,6,6,7,7,7,7,8,8,9,9,9,10,10,10,11,11,12,12,13,13,13,14,14,15,15,16,16),
            (7,7,6,6,6,6,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,14,14,15,15,16,16),
            (7,6,6,6,6,5,5,5,4,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,10,11,11,12,12,13,13,14,14,14,15,15,16),
            (7,6,6,6,5,5,5,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,12,13,13,14,14,15,15,16),
            (6,6,6,5,5,5,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6,7,7,8,8,8,9,9,10,10,10,11,11,12,12,13,13,14,14,15,15,16),
            (6,6,5,5,5,4,4,4,4,3,3,3,3,3,3,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,5,5,5,5,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,13,14,14,15,15),
            (6,5,5,5,4,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,10,10,11,11,11,12,12,13,13,14,14,15,15),
            (6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,14,14,15,15),
            (5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,2,2,2,1,1,1,2,2,2,2,2,2,2,3,3,3,3,4,4,4,4,5,5,6,6,6,7,7,8,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15,15),
            (5,5,5,4,4,4,3,3,3,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10,10,11,11,11,12,12,13,13,14,14,15),
            (5,5,4,4,4,3,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,5,5,5,6,6,6,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,4,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,3,3,3,3,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,0,0,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,4,3,3,3,2,2,2,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,3,3,3,3,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,12,13,13,14,15),
            (5,4,4,3,3,3,3,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,4,3,3,3,2,2,2,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,0,0,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,3,3,3,3,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,4,4,4,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,5,4,4,4,3,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,5,5,5,6,6,6,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,14,14,15),
            (5,5,5,4,4,4,3,3,3,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10,10,11,11,11,12,12,13,13,14,14,15),
            (5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,2,2,2,1,1,1,2,2,2,2,2,2,2,3,3,3,3,4,4,4,4,5,5,6,6,6,7,7,8,8,8,9,9,10,10,11,11,12,12,13,13,14,14,15,15),
            (6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,14,14,15,15),
            (6,5,5,5,4,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,10,10,11,11,11,12,12,13,13,14,14,15,15),
            (6,6,5,5,5,4,4,4,4,3,3,3,3,3,3,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,5,5,5,5,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,13,13,13,14,14,15,15),
            (6,6,6,5,5,5,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6,7,7,8,8,8,9,9,10,10,10,11,11,12,12,13,13,14,14,15,15,16),
            (7,6,6,6,5,5,5,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,9,9,9,10,10,11,11,12,12,12,13,13,14,14,15,15,16),
            (7,6,6,6,6,5,5,5,4,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,10,11,11,12,12,13,13,14,14,14,15,15,16),
            (7,7,6,6,6,6,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,14,14,15,15,16,16),
            (7,7,7,6,6,6,6,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,6,6,6,7,7,7,7,8,8,9,9,9,10,10,10,11,11,12,12,13,13,13,14,14,15,15,16,16),
            (8,7,7,7,6,6,6,6,5,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,10,10,10,11,11,12,12,12,13,13,14,14,15,15,16,16,16),
            (8,8,7,7,7,7,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,14,14,14,15,15,16,16,17),
            (8,8,8,7,7,7,7,6,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,11,11,11,12,12,13,13,13,14,14,15,15,16,16,16,17),
            (9,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,5,5,5,6,6,6,6,6,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,12,12,12,13,13,14,14,14,15,15,16,16,17,17),
            (9,9,8,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,8,8,8,9,9,9,9,10,10,10,11,11,12,12,12,13,13,13,14,14,15,15,16,16,17,17,17),
            (9,9,9,9,8,8,8,8,7,7,7,7,7,7,7,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,8,8,8,8,9,9,9,9,10,10,10,11,11,11,12,12,13,13,13,14,14,15,15,15,16,16,17,17,18),
            (10,9,9,9,9,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,9,9,9,10,10,10,10,11,11,11,12,12,13,13,13,14,14,14,15,15,16,16,17,17,17,18),
            (10,10,10,9,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,9,9,9,9,10,10,10,11,11,11,11,12,12,13,13,13,14,14,14,15,15,16,16,16,17,17,18,18),
            (10,10,10,10,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,10,10,10,10,11,11,11,12,12,12,13,13,13,14,14,14,15,15,16,16,16,17,17,18,18,18),
            (11,11,10,10,10,10,9,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,10,10,10,10,10,11,11,11,12,12,12,13,13,13,14,14,14,15,15,15,16,16,17,17,17,18,18,19),
            (11,11,11,11,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,11,11,11,11,12,12,12,13,13,13,14,14,14,15,15,15,16,16,17,17,17,18,18,19,19),
            (12,11,11,11,11,10,10,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,11,11,11,11,12,12,12,12,13,13,13,14,14,14,15,15,15,16,16,17,17,17,18,18,19,19,19),
            (12,12,12,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,9,9,9,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,12,12,12,12,13,13,13,14,14,14,15,15,15,16,16,16,17,17,18,18,18,19,19,20),
            (13,12,12,12,12,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,12,12,12,12,13,13,13,13,14,14,14,15,15,15,16,16,16,17,17,18,18,18,19,19,20,20),
            (13,13,12,12,12,12,12,11,11,11,11,11,11,11,11,11,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,12,12,12,12,12,13,13,13,13,14,14,14,14,15,15,15,16,16,16,17,17,18,18,18,19,19,20,20,20),
            (13,13,13,13,12,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,13,13,13,13,13,14,14,14,15,15,15,16,16,16,16,17,17,18,18,18,19,19,19,20,20,21),
            (14,14,13,13,13,13,13,12,12,12,12,12,12,12,12,12,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,13,13,13,13,13,14,14,14,14,15,15,15,16,16,16,17,17,17,18,18,18,19,19,19,20,20,21,21),
            (14,14,14,14,13,13,13,13,13,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,14,14,14,14,15,15,15,15,16,16,16,17,17,17,18,18,18,19,19,19,20,20,21,21,21),
            (15,14,14,14,14,14,14,13,13,13,13,13,13,13,13,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,14,14,14,14,14,15,15,15,15,16,16,16,16,17,17,17,18,18,18,19,19,19,20,20,21,21,21,22),
            (15,15,15,15,14,14,14,14,14,14,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,15,15,15,15,16,16,16,16,17,17,17,17,18,18,18,19,19,19,20,20,21,21,21,22,22),
            (16,15,15,15,15,15,14,14,14,14,14,14,14,14,14,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,16,16,16,16,17,17,17,18,18,18,19,19,19,19,20,20,21,21,21,22,22,22),
            (16,16,16,15,15,15,15,15,15,15,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,16,16,16,16,16,17,17,17,17,18,18,18,19,19,19,20,20,20,21,21,21,22,22,22,23));
            
     constant delay_matrix_3 : delay_matrix(0 to x_res-1) := ((24,23,23,22,22,22,21,21,21,20,20,20,19,19,19,18,18,18,18,17,17,17,17,16,16,16,16,16,15,15,15,15,15,15,15,15,15,15,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16),
            (23,23,22,22,22,21,21,21,20,20,20,19,19,19,18,18,18,17,17,17,17,16,16,16,16,16,15,15,15,15,15,15,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,16,16),
            (23,22,22,22,21,21,21,20,20,19,19,19,19,18,18,18,17,17,17,16,16,16,16,15,15,15,15,15,15,14,14,14,14,14,14,14,14,14,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,15,15,15,15,15),
            (22,22,22,21,21,21,20,20,19,19,19,18,18,18,17,17,17,17,16,16,16,16,15,15,15,15,14,14,14,14,14,14,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,15,15,15),
            (22,22,21,21,21,20,20,19,19,19,18,18,18,17,17,17,16,16,16,16,15,15,15,15,14,14,14,14,14,13,13,13,13,13,13,13,13,13,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,14,14,14,14,14,14),
            (22,21,21,21,20,20,19,19,19,18,18,18,17,17,17,16,16,16,15,15,15,15,14,14,14,14,13,13,13,13,13,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,14,14,14),
            (21,21,21,20,20,19,19,19,18,18,18,17,17,17,16,16,16,15,15,15,14,14,14,14,13,13,13,13,13,12,12,12,12,12,12,12,12,12,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,13,13,13,13,13,14),
            (21,21,20,20,19,19,19,18,18,18,17,17,16,16,16,16,15,15,15,14,14,14,13,13,13,13,13,12,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,13,13,13),
            (21,20,20,20,19,19,18,18,18,17,17,16,16,16,15,15,15,14,14,14,14,13,13,13,13,12,12,12,12,12,11,11,11,11,11,11,11,11,11,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,12,12,12,12,12,13),
            (20,20,20,19,19,18,18,18,17,17,16,16,16,15,15,15,14,14,14,13,13,13,13,12,12,12,12,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,12,12,12,12),
            (20,20,19,19,18,18,18,17,17,16,16,16,15,15,15,14,14,14,13,13,13,12,12,12,12,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,9,9,9,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,12,12),
            (20,19,19,19,18,18,17,17,17,16,16,15,15,15,14,14,14,13,13,13,12,12,12,12,11,11,11,11,10,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,11,11,11,11),
            (19,19,19,18,18,17,17,17,16,16,15,15,15,14,14,14,13,13,13,12,12,12,11,11,11,11,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,11,11,11),
            (19,19,18,18,17,17,17,16,16,15,15,15,14,14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,10,9,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,10,10,10,10,11),
            (19,18,18,18,17,17,16,16,16,15,15,14,14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,10,10,10),
            (19,18,18,17,17,16,16,16,15,15,14,14,14,13,13,13,12,12,11,11,11,11,10,10,10,9,9,9,9,8,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,9,9,9,9,10,10),
            (18,18,17,17,17,16,16,15,15,14,14,14,13,13,13,12,12,11,11,11,10,10,10,10,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,9,9,9,9),
            (18,18,17,17,16,16,15,15,15,14,14,13,13,13,12,12,11,11,11,10,10,10,9,9,9,9,8,8,8,8,7,7,7,7,7,7,7,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,8,8,8,8,9,9,9),
            (18,17,17,17,16,16,15,15,14,14,13,13,13,12,12,12,11,11,10,10,10,9,9,9,9,8,8,8,7,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,8,9),
            (18,17,17,16,16,15,15,14,14,14,13,13,12,12,12,11,11,10,10,10,9,9,9,8,8,8,8,7,7,7,7,6,6,6,6,6,6,6,6,6,5,5,5,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8),
            (17,17,16,16,16,15,15,14,14,13,13,13,12,12,11,11,11,10,10,9,9,9,8,8,8,8,7,7,7,7,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,7,7,7,7,8,8),
            (17,17,16,16,15,15,14,14,14,13,13,12,12,11,11,11,10,10,9,9,9,8,8,8,7,7,7,7,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8),
            (17,16,16,16,15,15,14,14,13,13,12,12,12,11,11,10,10,10,9,9,8,8,8,7,7,7,7,6,6,6,6,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,6,6,6,6,7,7,7),
            (17,16,16,15,15,14,14,13,13,13,12,12,11,11,10,10,10,9,9,9,8,8,7,7,7,7,6,6,6,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7),
            (17,16,16,15,15,14,14,13,13,12,12,11,11,11,10,10,9,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,6,6,6,6,7),
            (16,16,15,15,14,14,14,13,13,12,12,11,11,10,10,10,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,6,6,6,6),
            (16,16,15,15,14,14,13,13,12,12,12,11,11,10,10,9,9,9,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6),
            (16,16,15,15,14,14,13,13,12,12,11,11,10,10,10,9,9,8,8,8,7,7,6,6,6,5,5,5,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,6,6),
            (16,15,15,14,14,13,13,13,12,12,11,11,10,10,9,9,9,8,8,7,7,7,6,6,5,5,5,5,4,4,4,3,3,3,3,3,3,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,5,5,5,6),
            (16,15,15,14,14,13,13,12,12,11,11,11,10,10,9,9,8,8,7,7,7,6,6,6,5,5,5,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5),
            (16,15,15,14,14,13,13,12,12,11,11,10,10,9,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5),
            (16,15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,8,7,7,6,6,6,5,5,4,4,4,4,3,3,3,3,2,2,2,2,2,2,2,1,1,1,2,2,2,2,2,2,2,2,3,3,3,3,4,4,4,5,5),
            (15,15,14,14,13,13,12,12,11,11,11,10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,4,4,4,5,5),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,9,8,8,7,7,6,6,6,5,5,5,4,4,3,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,5),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,4,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,3,3,3,3,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,0,0,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,2,2,2,3,3,3,4,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,3,3,3,3,4,4),
            (15,15,14,13,13,12,12,12,11,11,10,10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,3,3,3,3,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,2,2,2,3,3,3,4,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,0,0,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,3,3,3,3,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,4,4,4),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5),
            (15,15,14,14,13,13,12,12,11,11,10,10,9,9,9,8,8,7,7,6,6,6,5,5,5,4,4,3,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,5),
            (15,15,14,14,13,13,12,12,11,11,11,10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,4,4,4,5,5),
            (16,15,15,14,14,13,13,12,12,11,11,10,10,9,9,8,8,8,7,7,6,6,6,5,5,4,4,4,4,3,3,3,3,2,2,2,2,2,2,2,1,1,1,2,2,2,2,2,2,2,2,3,3,3,3,4,4,4,5,5),
            (16,15,15,14,14,13,13,12,12,11,11,10,10,9,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5),
            (16,15,15,14,14,13,13,12,12,11,11,11,10,10,9,9,8,8,7,7,7,6,6,6,5,5,5,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5),
            (16,15,15,14,14,13,13,13,12,12,11,11,10,10,9,9,9,8,8,7,7,7,6,6,5,5,5,5,4,4,4,3,3,3,3,3,3,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,4,4,4,4,5,5,5,6),
            (16,16,15,15,14,14,13,13,12,12,11,11,10,10,10,9,9,8,8,8,7,7,6,6,6,5,5,5,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,6,6),
            (16,16,15,15,14,14,13,13,12,12,12,11,11,10,10,9,9,9,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6),
            (16,16,15,15,14,14,14,13,13,12,12,11,11,10,10,10,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,6,6,6,6),
            (17,16,16,15,15,14,14,13,13,12,12,11,11,11,10,10,9,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,6,6,6,6,7),
            (17,16,16,15,15,14,14,13,13,13,12,12,11,11,10,10,10,9,9,9,8,8,7,7,7,7,6,6,6,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7),
            (17,16,16,16,15,15,14,14,13,13,12,12,12,11,11,10,10,10,9,9,8,8,8,7,7,7,7,6,6,6,6,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,6,6,6,6,7,7,7),
            (17,17,16,16,15,15,14,14,14,13,13,12,12,11,11,11,10,10,9,9,9,8,8,8,7,7,7,7,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8),
            (17,17,16,16,16,15,15,14,14,13,13,13,12,12,11,11,11,10,10,9,9,9,8,8,8,8,7,7,7,7,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,7,7,7,7,8,8),
            (18,17,17,16,16,15,15,14,14,14,13,13,12,12,12,11,11,10,10,10,9,9,9,8,8,8,8,7,7,7,7,6,6,6,6,6,6,6,6,6,5,5,5,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8),
            (18,17,17,17,16,16,15,15,14,14,13,13,13,12,12,12,11,11,10,10,10,9,9,9,9,8,8,8,7,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,8,9),
            (18,18,17,17,16,16,15,15,15,14,14,13,13,13,12,12,11,11,11,10,10,10,9,9,9,9,8,8,8,8,7,7,7,7,7,7,7,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,8,8,8,8,9,9,9),
            (18,18,17,17,17,16,16,15,15,14,14,14,13,13,13,12,12,11,11,11,10,10,10,10,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,9,9,9,9),
            (19,18,18,17,17,16,16,16,15,15,14,14,14,13,13,13,12,12,11,11,11,11,10,10,10,9,9,9,9,8,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,9,9,9,9,10,10),
            (19,18,18,18,17,17,16,16,16,15,15,14,14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,10,10,10),
            (19,19,18,18,17,17,17,16,16,15,15,15,14,14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,10,9,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,10,10,10,10,11),
            (19,19,19,18,18,17,17,17,16,16,15,15,15,14,14,14,13,13,13,12,12,12,11,11,11,11,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,11,11,11),
            (20,19,19,19,18,18,17,17,17,16,16,15,15,15,14,14,14,13,13,13,12,12,12,12,11,11,11,11,10,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,11,11,11,11),
            (20,20,19,19,18,18,18,17,17,16,16,16,15,15,15,14,14,14,13,13,13,12,12,12,12,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,9,9,9,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,12,12),
            (20,20,20,19,19,18,18,18,17,17,16,16,16,15,15,15,14,14,14,13,13,13,13,12,12,12,12,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,12,12,12,12),
            (21,20,20,20,19,19,18,18,18,17,17,16,16,16,15,15,15,14,14,14,14,13,13,13,13,12,12,12,12,12,11,11,11,11,11,11,11,11,11,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,12,12,12,12,12,13),
            (21,21,20,20,19,19,19,18,18,18,17,17,16,16,16,16,15,15,15,14,14,14,13,13,13,13,13,12,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,13,13,13),
            (21,21,21,20,20,19,19,19,18,18,18,17,17,17,16,16,16,15,15,15,14,14,14,14,13,13,13,13,13,12,12,12,12,12,12,12,12,12,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,13,13,13,13,13,14),
            (22,21,21,21,20,20,19,19,19,18,18,18,17,17,17,16,16,16,15,15,15,15,14,14,14,14,13,13,13,13,13,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,14,14,14),
            (22,22,21,21,21,20,20,19,19,19,18,18,18,17,17,17,16,16,16,16,15,15,15,15,14,14,14,14,14,13,13,13,13,13,13,13,13,13,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,14,14,14,14,14,14),
            (22,22,22,21,21,21,20,20,19,19,19,18,18,18,17,17,17,17,16,16,16,16,15,15,15,15,14,14,14,14,14,14,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,15,15,15),
            (23,22,22,22,21,21,21,20,20,19,19,19,19,18,18,18,17,17,17,16,16,16,16,15,15,15,15,15,15,14,14,14,14,14,14,14,14,14,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,15,15,15,15,15),
            (23,23,22,22,22,21,21,21,20,20,20,19,19,19,18,18,18,17,17,17,17,16,16,16,16,16,15,15,15,15,15,15,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,16,16));
            
    constant delay_matrix_4 : delay_matrix(0 to x_res-1) := ((15,15,14,14,14,13,13,13,13,12,12,12,11,11,11,11,10,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,11,11,11,11,12,12,12,13,13,13,13,14,14,14,15),
            (15,14,14,14,13,13,13,12,12,12,12,11,11,11,10,10,10,10,10,9,9,9,9,9,9,9,9,9,8,8,8,8,8,9,9,9,9,9,9,9,9,9,10,10,10,10,10,11,11,11,12,12,12,12,13,13,13,14,14,14),
            (15,14,14,13,13,13,12,12,12,11,11,11,11,10,10,10,10,9,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,10,10,10,10,11,11,11,11,12,12,12,13,13,13,14,14),
            (14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,10,10,10,10,11,11,11,12,12,12,13,13,13,14),
            (14,13,13,13,12,12,12,11,11,11,10,10,10,10,9,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,9,9,9,9,10,10,10,10,11,11,11,12,12,12,13,13,13),
            (14,13,13,12,12,12,11,11,11,10,10,10,9,9,9,9,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,9,9,9,9,10,10,10,11,11,11,12,12,12,13,13),
            (13,13,12,12,12,11,11,11,10,10,10,9,9,9,8,8,8,8,8,7,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,8,8,8,8,8,9,9,9,10,10,10,11,11,11,12,12,12,13),
            (13,13,12,12,11,11,11,10,10,10,9,9,9,8,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,11,12,12,13),
            (13,12,12,11,11,11,10,10,10,9,9,9,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,5,5,5,5,5,5,5,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,11,12,12),
            (12,12,12,11,11,10,10,10,9,9,9,8,8,8,7,7,7,7,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,12,12),
            (12,12,11,11,10,10,10,9,9,9,8,8,8,7,7,7,7,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,10,11,11,12),
            (12,11,11,11,10,10,9,9,9,8,8,8,7,7,7,6,6,6,6,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,6,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11,11),
            (12,11,11,10,10,10,9,9,8,8,8,7,7,7,6,6,6,6,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,6,6,6,6,7,7,7,8,8,8,9,9,10,10,10,11,11),
            (11,11,11,10,10,9,9,9,8,8,7,7,7,6,6,6,6,5,5,5,5,4,4,4,4,4,4,4,4,3,3,3,4,4,4,4,4,4,4,4,5,5,5,5,6,6,6,6,7,7,7,8,8,9,9,9,10,10,11,11),
            (11,11,10,10,9,9,9,8,8,7,7,7,6,6,6,6,5,5,5,4,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,6,6,6,6,7,7,7,8,8,9,9,9,10,10,11),
            (11,10,10,10,9,9,8,8,8,7,7,7,6,6,6,5,5,5,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,10),
            (11,10,10,9,9,9,8,8,7,7,7,6,6,6,5,5,5,4,4,4,4,3,3,3,3,3,3,3,3,3,2,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,9,10,10),
            (11,10,10,9,9,8,8,8,7,7,6,6,6,5,5,5,4,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5,6,6,6,7,7,8,8,8,9,9,10,10),
            (10,10,9,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,9,10),
            (10,10,9,9,8,8,8,7,7,6,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,8,9,9,10),
            (10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,2,2,1,1,1,1,1,2,2,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10),
            (10,10,9,9,8,8,7,7,6,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,2,2,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,9,9,10),
            (10,9,9,8,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,8,9,9),
            (10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,3,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,3,4,4,5,5,5,6,6,7,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,0,0,0,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (9,9,9,8,8,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,9,9),
            (9,9,9,8,8,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,9,9),
            (9,9,9,8,8,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9),
            (10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9),
            (10,9,9,8,8,8,7,7,6,6,5,5,5,4,4,4,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,7,7,8,8,8,9,9),
            (10,9,9,9,8,8,7,7,6,6,6,5,5,4,4,4,3,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,5,5,6,6,6,7,7,8,8,9,9,9),
            (10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,2,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,4,4,4,5,5,5,6,6,7,7,7,8,8,9,9,10),
            (10,10,9,9,8,8,8,7,7,6,6,6,5,5,4,4,4,4,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,4,4,4,4,5,5,6,6,6,7,7,8,8,8,9,9,10),
            (10,10,9,9,9,8,8,7,7,6,6,6,5,5,5,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,9,9,9,10),
            (10,10,10,9,9,8,8,7,7,7,6,6,6,5,5,5,4,4,4,3,3,3,3,3,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,10,10),
            (11,10,10,9,9,8,8,8,7,7,7,6,6,5,5,5,5,4,4,4,3,3,3,3,3,3,3,2,2,2,2,2,2,2,3,3,3,3,3,3,3,4,4,4,5,5,5,5,6,6,7,7,7,8,8,8,9,9,10,10),
            (11,10,10,10,9,9,8,8,7,7,7,6,6,6,5,5,5,4,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,5,5,5,6,6,6,7,7,7,8,8,9,9,10,10,10),
            (11,11,10,10,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,11),
            (11,11,10,10,10,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,4,4,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,10,10,10,11),
            (11,11,11,10,10,9,9,9,8,8,8,7,7,7,6,6,6,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,6,6,6,7,7,7,8,8,8,9,9,9,10,10,11,11),
            (12,11,11,10,10,10,9,9,9,8,8,7,7,7,7,6,6,6,5,5,5,5,5,5,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,6,6,6,7,7,7,7,8,8,9,9,9,10,10,10,11,11),
            (12,12,11,11,10,10,10,9,9,8,8,8,7,7,7,7,6,6,6,6,5,5,5,5,5,5,5,4,4,4,4,4,4,4,5,5,5,5,5,5,5,6,6,6,6,7,7,7,7,8,8,8,9,9,10,10,10,11,11,12),
            (12,12,11,11,11,10,10,9,9,9,8,8,8,7,7,7,7,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,7,7,7,7,8,8,8,9,9,9,10,10,11,11,11,12),
            (12,12,12,11,11,11,10,10,9,9,9,8,8,8,8,7,7,7,7,6,6,6,6,6,6,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,7,7,7,7,8,8,8,8,9,9,9,10,10,11,11,11,12,12),
            (13,12,12,12,11,11,10,10,10,9,9,9,8,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,8,9,9,9,10,10,10,11,11,12,12,12),
            (13,13,12,12,12,11,11,10,10,10,9,9,9,9,8,8,8,8,7,7,7,7,7,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,8,8,8,8,9,9,9,9,10,10,10,11,11,12,12,12,13),
            (13,13,13,12,12,11,11,11,10,10,10,9,9,9,9,8,8,8,8,7,7,7,7,7,7,7,7,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,8,8,8,8,9,9,9,9,10,10,10,11,11,11,12,12,13,13),
            (14,13,13,13,12,12,11,11,11,10,10,10,10,9,9,9,9,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,9,9,9,9,10,10,10,10,11,11,11,12,12,13,13,13),
            (14,14,13,13,13,12,12,11,11,11,11,10,10,10,9,9,9,9,9,8,8,8,8,8,8,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,9,9,9,9,9,10,10,10,11,11,11,11,12,12,13,13,13,14),
            (14,14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,10,10,10,10,11,11,11,12,12,12,13,13,13,14,14),
            (15,14,14,14,13,13,13,12,12,12,11,11,11,10,10,10,10,10,9,9,9,9,9,9,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,10,10,10,10,10,11,11,11,12,12,12,13,13,13,14,14,14),
            (15,15,14,14,14,13,13,13,12,12,12,11,11,11,11,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,11,11,11,11,12,12,12,13,13,13,14,14,14,15),
            (15,15,15,14,14,14,13,13,13,12,12,12,12,11,11,11,11,10,10,10,10,10,10,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,11,11,11,11,12,12,12,12,13,13,13,14,14,14,15,15),
            (16,15,15,15,14,14,14,13,13,13,13,12,12,12,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,12,12,12,13,13,13,13,14,14,14,15,15,15),
            (16,16,15,15,15,14,14,14,13,13,13,13,12,12,12,12,12,11,11,11,11,11,11,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,12,12,12,12,12,13,13,13,13,14,14,14,15,15,15,16),
            (16,16,16,15,15,15,14,14,14,14,13,13,13,13,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,13,13,13,13,14,14,14,14,15,15,15,16,16),
            (17,17,16,16,16,15,15,15,14,14,14,14,13,13,13,13,12,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,13,13,13,13,14,14,14,14,15,15,15,16,16,16,17),
            (17,17,17,16,16,16,15,15,15,14,14,14,14,13,13,13,13,13,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,14,14,14,14,15,15,15,16,16,16,17,17),
            (18,17,17,17,16,16,16,15,15,15,15,14,14,14,14,14,13,13,13,13,13,13,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,14,14,14,14,14,15,15,15,15,16,16,16,17,17,17),
            (18,18,17,17,17,16,16,16,16,15,15,15,15,14,14,14,14,14,13,13,13,13,13,13,13,13,13,13,13,13,12,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,15,15,15,15,16,16,16,16,17,17,17,18),
            (18,18,18,17,17,17,17,16,16,16,16,15,15,15,15,14,14,14,14,14,14,14,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,15,15,15,15,16,16,16,16,17,17,17,17,18,18),
            (19,19,18,18,18,17,17,17,17,16,16,16,16,15,15,15,15,15,14,14,14,14,14,14,14,14,14,14,14,14,13,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,16,16,16,16,17,17,17,17,18,18,18,19),
            (19,19,19,18,18,18,17,17,17,17,16,16,16,16,16,15,15,15,15,15,15,15,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,16,16,16,16,16,17,17,17,17,18,18,18,19,19),
            (20,19,19,19,18,18,18,18,17,17,17,17,16,16,16,16,16,16,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,17,17,17,17,18,18,18,18,19,19,19),
            (20,20,19,19,19,19,18,18,18,18,17,17,17,17,17,16,16,16,16,16,16,16,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,17,17,17,17,17,18,18,18,18,19,19,19,19,20),
            (21,20,20,20,19,19,19,19,18,18,18,18,17,17,17,17,17,17,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,17,17,17,17,17,18,18,18,18,19,19,19,19,20,20,20),
            (21,21,20,20,20,20,19,19,19,19,18,18,18,18,18,17,17,17,17,17,17,17,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,17,17,17,17,17,17,18,18,18,18,18,19,19,19,19,20,20,20,20,21),
            (21,21,21,21,20,20,20,20,19,19,19,19,18,18,18,18,18,18,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,18,18,18,18,18,18,19,19,19,19,20,20,20,20,21,21,21),
            (22,22,21,21,21,20,20,20,20,20,19,19,19,19,19,18,18,18,18,18,18,18,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,18,18,18,18,18,18,18,19,19,19,19,19,20,20,20,20,20,21,21,21,22),
            (22,22,22,21,21,21,21,20,20,20,20,20,19,19,19,19,19,19,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,19,19,19,19,19,19,20,20,20,20,20,21,21,21,21,22,22),
            (23,22,22,22,22,21,21,21,21,20,20,20,20,20,20,19,19,19,19,19,19,19,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,19,19,19,19,19,19,19,20,20,20,20,20,20,21,21,21,21,22,22,22,22),
            (23,23,23,22,22,22,22,21,21,21,21,21,20,20,20,20,20,20,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,20,20,20,20,20,20,21,21,21,21,21,22,22,22,22,23,23),
            (24,23,23,23,23,22,22,22,22,21,21,21,21,21,21,20,20,20,20,20,20,20,20,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,20,20,20,20,20,20,20,20,21,21,21,21,21,21,22,22,22,22,23,23,23,23),
            (24,24,24,23,23,23,23,22,22,22,22,22,21,21,21,21,21,21,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,21,21,21,21,21,22,22,22,22,22,23,23,23,23,24,24));

    constant max_delay : integer := 25;
    
    type input_buffer_array is array (0 to max_delay) of signed(15 downto 0);
                 
end package;

package body pkg is
end package body;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

library work;
use work.pkg.all;


entity beam_gen is
    Generic (   HEIGHT  :       INTEGER := 480;     -- screen hight
                WIDTH   :       INTEGER := 640;     -- screen width
                MAX_SEL :       integer := 0);
    Port ( clk_d :  in STD_LOGIC;
           clk_p :  in STD_LOGIC;
           nrst :   in STD_LOGIC;
           sound1 : in std_logic_vector(15 downto 0);
           sound2 : in std_logic_vector(15 downto 0);
           sound3 : in std_logic_vector(15 downto 0);
           sound4 : in std_logic_vector(15 downto 0);
           row :    in unsigned (9 downto 0);
           col :    in unsigned (9 downto 0);
           video:   out std_logic_vector(11 downto 0);
           nsample: in std_logic;
           disp_en: in std_logic;
           D_out :  out std_logic_vector(31 downto 0);
           sel :    in std_logic);
end beam_gen;

architecture Behavioral of beam_gen is
    
    signal input_buffer_1 : input_buffer_array  := (others => (others => '0'));
    signal input_buffer_2 : input_buffer_array  := (others => (others => '0'));
    signal input_buffer_3 : input_buffer_array  := (others => (others => '0'));
    signal input_buffer_4 : input_buffer_array  := (others => (others => '0'));
    
    signal signal_buffer_1 : input_buffer_array := (others => (others => '0'));
    signal signal_buffer_2 : input_buffer_array := (others => (others => '0'));
    signal signal_buffer_3 : input_buffer_array := (others => (others => '0'));
    signal signal_buffer_4 : input_buffer_array := (others => (others => '0'));
    
    signal sound_sum :      signed(15 downto 0) := (others => '0');
    
    signal output_buffer :  signed(31 downto 0) := (others => '0');
    
    signal ind_x :          unsigned(9 downto 0)    := (others => '0');
    signal ind_y :          unsigned(9 downto 0)    := (others => '0');
    
    signal const_buff_1 :   delay_array(0 to y_res-1);
    signal const_buff_2 :   delay_array(0 to y_res-1);
    signal const_buff_3 :   delay_array(0 to y_res-1);
    signal const_buff_4 :   delay_array(0 to y_res-1);
    
--    signal en :             std_logic               := '0';
    
    signal test_input_buffer : input_buffer_array  := (x"0fff",
                                                        x"0ff0",
                                                        x"0f00",
                                                        x"0e00",
                                                        x"0d00",
                                                        x"0c00",
                                                        x"0b00",
                                                        x"0a00",
                                                        x"0900",
                                                        x"0800",
                                                        x"00f0",
                                                        x"00e0",
                                                        x"00d0",
                                                        x"00c0",
                                                        x"00b0",
                                                        x"00a0",
                                                        x"0090",
                                                        x"0080",
                                                        x"000f",
                                                        x"000e",
                                                        x"000d",
                                                        x"000c",
                                                        x"000b",
                                                        x"000a",
                                                        x"0009",
                                                        x"0008");
    
begin

    ind_x <= b"000" & col(9 downto 3);
    ind_y <= b"000" & row(9 downto 3);
    
--buffering_ctrl: process(nsample, nrst)
--begin
--    if (nrst = '0') then
--        en <= '0';
--    elsif (nsample = '0') then
--        en <= '1';
--    else
--        en <= '0';
--    end if;
--end process;
    
input_buffering: process(clk_d, nrst)
begin 
    if (nrst = '0') then
    
        input_buffer_1 <= (others => (others => '0'));
        input_buffer_2 <= (others => (others => '0'));
        input_buffer_3 <= (others => (others => '0'));
        input_buffer_4 <= (others => (others => '0'));
        
    elsif (rising_edge(clk_d)) then
    
        if (nsample = '0') then
        
            for ii in 1 to max_delay loop
                input_buffer_1(ii) <= input_buffer_1(ii-1);
                input_buffer_2(ii) <= input_buffer_2(ii-1);
                input_buffer_3(ii) <= input_buffer_3(ii-1);
                input_buffer_4(ii) <= input_buffer_4(ii-1);
            end loop;
            
            input_buffer_1(0) <= signed(sound1);
            input_buffer_2(0) <= signed(sound2);
            input_buffer_3(0) <= signed(sound3);
            input_buffer_4(0) <= signed(sound4);
            
        end if;
    end if;
    
end process;

    const_buff_1 <= delay_matrix_1(to_integer(ind_x));
   --const_buff_1 <= delay_matrix_1(53);
    const_buff_2 <= delay_matrix_2(to_integer(ind_x));
    const_buff_3 <= delay_matrix_3(to_integer(ind_x));
    const_buff_4 <= delay_matrix_4(to_integer(ind_x));

delay_and_sum: process(clk_p, nrst)
begin 
    if (nrst = '0') then
    
        sound_sum <= (others => '0');
        
        signal_buffer_1 <= (others => (others => '0'));
        signal_buffer_2 <= (others => (others => '0'));
        signal_buffer_3 <= (others => (others => '0'));
        signal_buffer_4 <= (others => (others => '0'));
        
    elsif (rising_edge(clk_p)) then
    
        if (disp_en = '1') then
            if (to_integer(row) < (WIDTH)) then
        --sound_sum <= test_input_buffer(const_buff_1(50));                         -- this part works
                
                if ((row = to_unsigned(0, 10)) and (col = to_unsigned(0, 10))) then
                    signal_buffer_1 <= input_buffer_1;
                    signal_buffer_2 <= input_buffer_2;
                    signal_buffer_3 <= input_buffer_3;
                    signal_buffer_4 <= input_buffer_4;
                    
                end if;
                
                if (to_integer(ind_y) < HEIGHT) then
                    --sound_sum <= test_input_buffer(const_buff_3(to_integer(ind_y)));
                    --sound_sum <= x"ff0f";
--                    sound_sum <= test_input_buffer(const_buff_1(to_integer(ind_y))) +
--                        test_input_buffer(const_buff_2(to_integer(ind_y))) +
--                        test_input_buffer(const_buff_3(to_integer(ind_y))) +
--                        test_input_buffer(const_buff_4(to_integer(ind_y)));
                    sound_sum <= signal_buffer_1(const_buff_1(to_integer(ind_y))) +
                        signal_buffer_2(const_buff_2(to_integer(ind_y))) +
                        signal_buffer_3(const_buff_3(to_integer(ind_y))) +
                        signal_buffer_4(const_buff_4(to_integer(ind_y)));
                        
                 else
                    sound_sum <= x"0000";
                 end if;
            --sound_sum <= x"ffff";--test_input_buffer(0);
           --sound_sum <= test_input_buffer(const_buff_1(to_integer(ind_y))); --+
    --                input_buffer_2(const_buff_1(to_integer(ind_y))) +
    --                input_buffer_3(const_buff_1(to_integer(ind_y))) +
    --                input_buffer_4(const_buff_1(to_integer(ind_y)));
    --        sound_sum <= to_signed(const_buff_1(to_integer(ind_y)), 16) +
    --                to_signed(const_buff_2(to_integer(ind_y)), 16) +
    --                to_signed(const_buff_3(to_integer(ind_y)), 16) +
    --                to_signed(const_buff_4(to_integer(ind_y)), 16);
            else
                sound_sum <= x"0000";
            end if;
        else
            sound_sum <= x"0000";
        end if;
    end if;
end process;

    output_buffer <= sound_sum*sound_sum;
    
    with sel select
        video <= std_logic_vector(output_buffer(MAX_SEL+10+13 downto MAX_SEL+10+10)) & 
                std_logic_vector(output_buffer(MAX_SEL+10+9 downto MAX_SEL+10+6)) & 
                std_logic_vector(output_buffer(MAX_SEL+10+3 downto MAX_SEL+10)) when '1',
                std_logic_vector(output_buffer(MAX_SEL+15 downto MAX_SEL+12)) & 
                std_logic_vector(output_buffer(MAX_SEL+9 downto MAX_SEL+6)) & 
                std_logic_vector(output_buffer(MAX_SEL+3 downto MAX_SEL)) when '0',
                (others => '0') when others;
    --video <= std_logic_vector(output_buffer(MAX_SEL+11 downto MAX_SEL));
    --video <= std_logic_vector(sound_sum(MAX_SEL+11 downto MAX_SEL));
    
    D_out <= std_logic_vector(output_buffer);

end Behavioral;
